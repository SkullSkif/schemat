library verilog;
use verilog.vl_types.all;
entity mem32_t is
end mem32_t;
